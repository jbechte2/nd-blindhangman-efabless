magic
tech gf180mcuD
magscale 1 5
timestamp 1702320099
<< obsm1 >>
rect 672 1538 279328 174078
<< metal2 >>
rect 69888 0 69944 400
rect 209888 0 209944 400
<< obsm2 >>
rect 854 430 279146 174067
rect 854 400 69858 430
rect 69974 400 209858 430
rect 209974 400 279146 430
<< metal3 >>
rect 279600 171472 280000 171528
rect 279600 163520 280000 163576
rect 279600 155568 280000 155624
rect 0 154000 400 154056
rect 279600 147616 280000 147672
rect 279600 139664 280000 139720
rect 279600 131712 280000 131768
rect 279600 123760 280000 123816
rect 279600 115808 280000 115864
rect 0 109984 400 110040
rect 279600 107856 280000 107912
rect 279600 99904 280000 99960
rect 279600 91952 280000 92008
rect 279600 84000 280000 84056
rect 279600 76048 280000 76104
rect 279600 68096 280000 68152
rect 0 65968 400 66024
rect 279600 60144 280000 60200
rect 279600 52192 280000 52248
rect 279600 44240 280000 44296
rect 279600 36288 280000 36344
rect 279600 28336 280000 28392
rect 0 21952 400 22008
rect 279600 20384 280000 20440
rect 279600 12432 280000 12488
rect 279600 4480 280000 4536
<< obsm3 >>
rect 400 171558 279650 174062
rect 400 171442 279570 171558
rect 400 163606 279650 171442
rect 400 163490 279570 163606
rect 400 155654 279650 163490
rect 400 155538 279570 155654
rect 400 154086 279650 155538
rect 430 153970 279650 154086
rect 400 147702 279650 153970
rect 400 147586 279570 147702
rect 400 139750 279650 147586
rect 400 139634 279570 139750
rect 400 131798 279650 139634
rect 400 131682 279570 131798
rect 400 123846 279650 131682
rect 400 123730 279570 123846
rect 400 115894 279650 123730
rect 400 115778 279570 115894
rect 400 110070 279650 115778
rect 430 109954 279650 110070
rect 400 107942 279650 109954
rect 400 107826 279570 107942
rect 400 99990 279650 107826
rect 400 99874 279570 99990
rect 400 92038 279650 99874
rect 400 91922 279570 92038
rect 400 84086 279650 91922
rect 400 83970 279570 84086
rect 400 76134 279650 83970
rect 400 76018 279570 76134
rect 400 68182 279650 76018
rect 400 68066 279570 68182
rect 400 66054 279650 68066
rect 430 65938 279650 66054
rect 400 60230 279650 65938
rect 400 60114 279570 60230
rect 400 52278 279650 60114
rect 400 52162 279570 52278
rect 400 44326 279650 52162
rect 400 44210 279570 44326
rect 400 36374 279650 44210
rect 400 36258 279570 36374
rect 400 28422 279650 36258
rect 400 28306 279570 28422
rect 400 22038 279650 28306
rect 430 21922 279650 22038
rect 400 20470 279650 21922
rect 400 20354 279570 20470
rect 400 12518 279650 20354
rect 400 12402 279570 12518
rect 400 4566 279650 12402
rect 400 4450 279570 4566
rect 400 1554 279650 4450
<< metal4 >>
rect 2224 1538 2384 174078
rect 9904 1538 10064 174078
rect 17584 1538 17744 174078
rect 25264 1538 25424 174078
rect 32944 1538 33104 174078
rect 40624 1538 40784 174078
rect 48304 1538 48464 174078
rect 55984 1538 56144 174078
rect 63664 1538 63824 174078
rect 71344 1538 71504 174078
rect 79024 1538 79184 174078
rect 86704 1538 86864 174078
rect 94384 1538 94544 174078
rect 102064 1538 102224 174078
rect 109744 1538 109904 174078
rect 117424 1538 117584 174078
rect 125104 1538 125264 174078
rect 132784 1538 132944 174078
rect 140464 1538 140624 174078
rect 148144 1538 148304 174078
rect 155824 1538 155984 174078
rect 163504 1538 163664 174078
rect 171184 1538 171344 174078
rect 178864 1538 179024 174078
rect 186544 1538 186704 174078
rect 194224 1538 194384 174078
rect 201904 1538 202064 174078
rect 209584 1538 209744 174078
rect 217264 1538 217424 174078
rect 224944 1538 225104 174078
rect 232624 1538 232784 174078
rect 240304 1538 240464 174078
rect 247984 1538 248144 174078
rect 255664 1538 255824 174078
rect 263344 1538 263504 174078
rect 271024 1538 271184 174078
rect 278704 1538 278864 174078
<< obsm4 >>
rect 248934 68833 255634 84047
rect 255854 68833 263314 84047
rect 263534 68833 265202 84047
<< labels >>
rlabel metal3 s 279600 4480 280000 4536 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 65968 400 66024 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 21952 400 22008 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 279600 28336 280000 28392 6 io_in[1]
port 4 nsew signal input
rlabel metal3 s 279600 52192 280000 52248 6 io_in[2]
port 5 nsew signal input
rlabel metal3 s 279600 76048 280000 76104 6 io_in[3]
port 6 nsew signal input
rlabel metal3 s 279600 99904 280000 99960 6 io_in[4]
port 7 nsew signal input
rlabel metal3 s 279600 123760 280000 123816 6 io_in[5]
port 8 nsew signal input
rlabel metal3 s 279600 147616 280000 147672 6 io_in[6]
port 9 nsew signal input
rlabel metal3 s 279600 171472 280000 171528 6 io_in[7]
port 10 nsew signal input
rlabel metal3 s 0 154000 400 154056 6 io_in[8]
port 11 nsew signal input
rlabel metal3 s 0 109984 400 110040 6 io_in[9]
port 12 nsew signal input
rlabel metal3 s 279600 20384 280000 20440 6 io_oeb[0]
port 13 nsew signal output
rlabel metal3 s 279600 44240 280000 44296 6 io_oeb[1]
port 14 nsew signal output
rlabel metal3 s 279600 68096 280000 68152 6 io_oeb[2]
port 15 nsew signal output
rlabel metal3 s 279600 91952 280000 92008 6 io_oeb[3]
port 16 nsew signal output
rlabel metal3 s 279600 115808 280000 115864 6 io_oeb[4]
port 17 nsew signal output
rlabel metal3 s 279600 139664 280000 139720 6 io_oeb[5]
port 18 nsew signal output
rlabel metal3 s 279600 163520 280000 163576 6 io_oeb[6]
port 19 nsew signal output
rlabel metal3 s 279600 12432 280000 12488 6 io_out[0]
port 20 nsew signal output
rlabel metal3 s 279600 36288 280000 36344 6 io_out[1]
port 21 nsew signal output
rlabel metal3 s 279600 60144 280000 60200 6 io_out[2]
port 22 nsew signal output
rlabel metal3 s 279600 84000 280000 84056 6 io_out[3]
port 23 nsew signal output
rlabel metal3 s 279600 107856 280000 107912 6 io_out[4]
port 24 nsew signal output
rlabel metal3 s 279600 131712 280000 131768 6 io_out[5]
port 25 nsew signal output
rlabel metal3 s 279600 155568 280000 155624 6 io_out[6]
port 26 nsew signal output
rlabel metal4 s 2224 1538 2384 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 174078 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 174078 6 vss
port 28 nsew ground bidirectional
rlabel metal2 s 69888 0 69944 400 6 wb_clk_i
port 29 nsew signal input
rlabel metal2 s 209888 0 209944 400 6 wb_rst_i
port 30 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 280000 176000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16339414
string GDS_FILE /home/jbech002/nd-blindhangman-efabless/openlane/user_proj_example/runs/23_12_11_13_36/results/signoff/user_proj_example.magic.gds
string GDS_START 336912
<< end >>

